class apb_sequence extends uvm_sequence #(apb_seq_item);
  
  `uvm_object_utils(apb_sequence)
  
  function new(string name="apb_sequence");
    super.new(name);
  endfunction
  
   task body();
     repeat(500) begin
     req = apb_seq_item::type_id::create("req");
     start_item(req);
       assert(req.randomize());
     finish_item(req);
       //req.print();
     end

     
   endtask
    
    
endclass